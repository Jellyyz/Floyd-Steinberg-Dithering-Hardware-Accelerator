// `timescale 10ns/1ns
// module pixel_tb(); 
    
// pixel_algorithm_unit p0(
//     // input 
//     .clk(clk), .rst(rst), // clk-rst itf 
//     .color(color), 
//     // ouput 
//     .color(color_out)
// ); 

// task reset(); 
// 	forever begin 
// 		 #1 clk = ~clk; 
// 	end 

//     clk = 1'b0; 
//     rst = 1'b0; 
// #1  rst = 1'b1;
// #1  rst = 1'b0; 

// endtask

// task int_mem(); 
//     $display("Loading memory chunks..."); 
    
    
// endtask

// task mosi(); 

// endtask

// task miso(); 

// endtask


// initial begin: 

//     reset(); 
    
// #5  int_mem(); 






// end 




// endmodule 