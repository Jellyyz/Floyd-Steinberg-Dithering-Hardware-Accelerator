module mem_itf(
    input logic clk, rst,
    input logic mem_data_in, 
    input logic me


)