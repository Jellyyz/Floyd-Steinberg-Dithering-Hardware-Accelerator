module top(
    // CLk - Rst Interface 
    input logic CLk, Rst 
    input logic [7:0] red, green, blue 

); 

logic [31:0] png_data []

// reading stuff from a file section of code



endmodule 